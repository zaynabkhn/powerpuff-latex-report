module not_1b (
    input wire a,
    output wire y
);
    assign y = ~a;
endmodule
